`timescale 1ns/1ps

// SRI HARI A S

module otsu_tb();
    logic clk;
    logic rst_n;
    logic start;
    logic [7:0] pixel_in;
    logic pixel_valid;
    logic last_pixel;

    logic [7:0] threshold;
    logic done;

    localparam IMG_WIDTH  = 512;
    localparam IMG_HEIGHT = 512;
    localparam TOTAL_PIXELS = IMG_WIDTH * IMG_HEIGHT;

    logic [7:0] img_mem [0:TOTAL_PIXELS-1];

    otsu_thresholding_fpga dut (.*);

    initial clk = 0;
    always #5 clk = ~clk;

    initial begin
        rst_n = 0;
        start = 0;
        pixel_in = 0;
        pixel_valid = 0;
        last_pixel = 0;

        // Loading hex file (generated by Python)
        $readmemh("image_in.hex", img_mem);

        repeat(5) @(posedge clk);
        rst_n = 1;
        repeat(5) @(posedge clk);

        start = 1;
        @(posedge clk);
        start = 0;

        // Wait for CLEAR state to finish (256 cycles)
        wait(dut.state == dut.BUILD);

        $display("[%0t] Streaming %0d pixels...", $time, TOTAL_PIXELS);
        for (int i = 0; i < TOTAL_PIXELS; i++) begin
            @(posedge clk);
            pixel_in    <= img_mem[i];
            pixel_valid <= 1;
            if (i == TOTAL_PIXELS - 1)
                last_pixel <= 1;
        end

        @(posedge clk);
        pixel_valid <= 0;
        last_pixel  <= 0;

        wait(done);
        $display("--------------------------------------");
        $display("Hardware Threshold Found: %d", threshold);
        $display("--------------------------------------");
        
        repeat(10) @(posedge clk);
        $finish;
    end

endmodule
